module main(
    input logic [9:0] switches,
    input logic clkButton, PKb // reset button?
    output logic [9:0] leds,
    output logic [6:0] hexes [2:0], // 3 hex displays
    output logic [6:0] timeStepHex,
    output logic doneSignalDP
);


endmodule